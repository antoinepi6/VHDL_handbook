-- File: counter_arch.vhd

